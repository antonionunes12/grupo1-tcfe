Circuito L2 - Alterado
*
* NGSPICE simulation script
* Req Calculator
*

.options savecurrents

*Indepedent Voltage Source
Va 1 0 0
Vx 6 9 8.801255

*Resistors
R1 1 2 1.03504497262k
R2 3 2 2.01159104669k 
R3 2 5 3.03557466091k
R4 5 0 4.10235086526k
R5 5 6 3.09889833746k
R6 0 7 2.00952426524k
R7 8 9 1.04158528578k

*Dummy 0V-Voltage Source to Measure Current through R6 (Ic)
Vaux 7 8 0.0

*Current Controlled Voltage Source
Hc 5 9 Vaux 8.09359354837k

*Voltage Controlled Current Source
Gb 6 3 (2,5) 7.3172497028m


.model linearcircuit NPN
.control
op

echo "********************************************"
echo  "Operating point"
echo "********************************************"

echo "op_TAB"
print all
echo "op_END"
quit
.endc

.end
